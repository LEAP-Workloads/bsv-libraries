
interface PLB_DEVICE;
  interface PLBMasterWires plbMasterWires;
  interface PLBSlaveWires#(32,64) plbSlaveWires;  
endinterface
